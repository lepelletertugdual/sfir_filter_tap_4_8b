-- #################################################################################################################################################################################
-- file :
--     gen_heartbeat.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     indicates FPGA activity.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     register tranfer level (RTL)
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     clock ratio must be higher or equal to 16.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2023-11-11
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--     02. entity
--     03. architecture
--         03.01. constants
--         03.02. signals
--         03.03. input assignment
--         03.04. alive output pin generation
--         03.05. output assignment
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;

    -- =============================================================================================================================================================================
	-- 01.01. custom
    -- =============================================================================================================================================================================	
	library work;
	    use work.pkg_gen_heartbeat.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity gen_heartbeat is
    generic (
	     g_clk_i_freq : integer := 100_000_000
		;g_clk_o_freq : integer :=   5_000_000
	);
    port (
	     i_clk   : in  std_logic
		;i_rst   : in  std_logic
		;o_alive : out std_logic
		;o_error : out std_logic_vector(7 downto 0)
	);
end entity gen_heartbeat;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture rtl of gen_heartbeat is

    -- =============================================================================================================================================================================
	-- 03.01. constants
    -- =============================================================================================================================================================================
	constant c_clk_ratio : integer := integer(real(g_clk_i_freq)/real(g_clk_o_freq));

    -- =============================================================================================================================================================================
	-- 03.02. signals
    -- =============================================================================================================================================================================
	signal s_clk         : std_logic;
	signal s_rst         : std_logic;
    signal s_cnt         : integer range 0 to c_clk_ratio/2-1;
	signal s_alive       : std_logic;
	signal s_error_ratio : std_logic;

begin

    -- =============================================================================================================================================================================
	-- 03.03. check input parameters
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. check clock ratio
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    check_clk_ratio_ok : if (c_clk_ratio > c_clk_ratio_upper_bound or c_clk_ratio = c_clk_ratio_upper_bound) generate
	        s_error_ratio <= '0';
	    end generate check_clk_ratio_ok;

	    check_clk_ratio_ko : if (c_clk_ratio < c_clk_ratio_upper_bound) generate
	        s_error_ratio <= '1';
	    end generate check_clk_ratio_ko;

    -- =============================================================================================================================================================================
	-- 03.04. input assignment
    -- =============================================================================================================================================================================
	s_clk <= i_clk;
	s_rst <= i_rst;

    -- =============================================================================================================================================================================
	-- 03.05. alive output pin generation
    -- =============================================================================================================================================================================
    p_gen_alive : process(s_rst,s_clk)
	begin
	    if (s_rst = '1') then
		    s_cnt <= 0;
			s_alive <= '0';
		elsif (rising_edge(s_clk)) then
		    if (s_cnt = c_clk_ratio/2-1) then
			    s_cnt <= 0;
				s_alive <= not(s_alive);
			else
			    s_cnt <= s_cnt + 1;
			end if;
		end if;
	end process p_gen_alive;

    -- =============================================================================================================================================================================
	-- 03.06. output assignment
    -- =============================================================================================================================================================================
	o_alive <= s_alive;
    o_error <= (
	     c_pos_error_ratio => s_error_ratio
		,others            => '0'
	);

end architecture rtl;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################