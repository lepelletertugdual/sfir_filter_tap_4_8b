-- ######################################################################################################################################################################################################
-- file :
--     pkg_mgt_file.vhd
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     procedures definition for file management.
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     none
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     none
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2023-11-11
--         file creation
-- ------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--         01.01. standard
--     02. package header
--         02.01. procedure prototypes
--             02.01.01. LOG
--                 02.01.01.01. file_log_open
--                 02.01.01.02. file_log_close
--             02.02.01. RPT
--                 02.02.01.01. file_rpt_open
--                 02.02.01.02. file_rpt_close
--     03. package body
--         03.01. procedure definition
--             03.01.01. LOG
--                 03.01.01.01. file_log_open
--                 03.01.01.02. file_log_close
--             03.01.02. RPT
--                 03.01.02.01. file_rpt_open
--                 03.01.02.02. file_rpt_close
-- ######################################################################################################################################################################################################

-- ######################################################################################################################################################################################################
-- 01. libraries
-- ######################################################################################################################################################################################################
    -- ==================================================================================================================================================================================================
	-- 01.01. standard
    -- ==================================================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
        use ieee.numeric_std.all;

    library std;
        use std.textio.all;

-- ######################################################################################################################################################################################################
-- 02. package header
-- ######################################################################################################################################################################################################

package pkg_mgt_file is
    
    -- ==================================================================================================================================================================================================
	-- 02.01. procedure prototypes
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 02.01.01. LOG
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
            -- ==========================================================================================================================================================================================
	        -- 02.01.01.01. proc_file_log_open
            -- ==========================================================================================================================================================================================
            procedure proc_file_log_open (
                 constant c_file_name : string
		        ;file     f_file      : text
            );
    
            -- ==========================================================================================================================================================================================
	        -- 02.01.01.01. proc_file_log_close
            -- ==========================================================================================================================================================================================
            procedure proc_file_log_close (
                 constant c_file_name : string
		        ;file     f_file      : text
            );
    
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 02.01.02. RPT
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
            -- ==========================================================================================================================================================================================
	        -- 02.01.02.01. proc_file_rpt_open
            -- ==========================================================================================================================================================================================
            procedure proc_file_rpt_open (
                 constant c_file_name : string
		        ;file     f_file      : text
            );
    
            -- ==========================================================================================================================================================================================
	        -- 02.01.02.02. proc_file_rpt_close
            -- ==========================================================================================================================================================================================
            procedure proc_file_rpt_close (
                 constant c_file_name : string
		        ;file     f_file      : text
            );
	
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 02.01.02. STM
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
            -- ==========================================================================================================================================================================================
	        -- 02.01.02.01. proc_file_stm_open
            -- ==========================================================================================================================================================================================
            procedure proc_file_stm_open (
                 constant c_file_name : string
		        ;file     f_file      : text
            );
    
            -- ==========================================================================================================================================================================================
	        -- 02.01.02.02. proc_file_stm_close
            -- ==========================================================================================================================================================================================
            procedure proc_file_stm_close (
                 constant c_file_name : string
		        ;file     f_file      : text
            );
	
end package pkg_mgt_file;

-- ######################################################################################################################################################################################################
-- 03. package body
-- ######################################################################################################################################################################################################

package body pkg_mgt_file is

    -- ==================================================================================================================================================================================================
	-- 03.01. procedure definition
    -- ==================================================================================================================================================================================================
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. LOG
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
            -- ==========================================================================================================================================================================================
	        -- 03.01.01.01. proc_file_log_open
            -- ==========================================================================================================================================================================================
            procedure proc_file_log_open (
                 constant c_file_name : string
		        ;file     f_file      : text
            ) is                  
			    constant c_field_separator : string := " ";
				constant c_proc_name       : string := "proc_file_log_open";
                variable v_file_status     : file_open_status;
            begin
                file_open(v_file_status,f_file,c_file_name,write_mode);
		        -- successfully opened
                if (v_file_status = OPEN_OK) then
                    assert false
			            report c_file_name                   & -- file name 
						           c_field_separator         & -- field separator
							           c_proc_name           & -- procedure name
									       c_field_separator & -- field separator
										       "success"       -- message
				        severity note;
                -- error
                else
		            -- status error
                    if (v_file_status = STATUS_ERROR) then
                        assert false
			                report c_file_name                              & -- file name
							           c_field_separator                    & -- field separator
									       c_proc_name                      & -- procedure name
										       c_field_separator            & -- field separator
											       "failure : status_error"   -- message
				            severity failure;
                    -- name error 
                    elsif (v_file_status = NAME_ERROR) then
                        assert false
			                report c_file_name                              & -- file name
							           c_field_separator                    & -- field separator
									       c_proc_name                      & -- procedure name
										       c_field_separator            & -- field separator
											       "failure : name_error"     -- message
				                severity failure;
			        -- failed to open
                    else
                        assert false
			                report c_file_name                   & -- file name
 							           c_field_separator         & -- field separator 
									       c_proc_name           & -- procedure name
										       c_field_separator & -- field separator
 											       "failure"       -- message
				            severity failure;
                    end if;
		        end if;
            end procedure proc_file_log_open;

            -- ==========================================================================================================================================================================================
	        -- 03.01.01.02. proc_file_log_close
            -- ==========================================================================================================================================================================================
            procedure proc_file_log_close (
                 constant c_file_name : string
		        ;file     f_file      : text
            ) is 
				constant c_proc_name       : string := "proc_file_log_close";
			    constant c_field_separator : string := " ";			
            begin
                file_close(f_file);
		        assert false
			        report c_file_name                   & -- file name
                               c_field_separator         & -- field separator
							       c_proc_name           & -- procedure name
								       c_field_separator & -- field separator
									       "success"       -- message
			        severity note;
            end procedure proc_file_log_close;
    
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.02. RPT
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
            -- ==========================================================================================================================================================================================
	        -- 03.01.02.01. proc_file_rpt_open
            -- ==========================================================================================================================================================================================
            procedure proc_file_rpt_open (
                 constant c_file_name : string
		        ;file     f_file      : text
            ) is                  
				constant c_proc_name       : string := "proc_file_rpt_open";
			    constant c_field_separator : string := " ";
                variable v_file_status     : file_open_status;
            begin
                file_open(v_file_status,f_file,c_file_name,write_mode);
		        -- successfully opened
                if (v_file_status = OPEN_OK) then
                    assert false
			            report c_file_name                   & -- file name 
						           c_field_separator         & -- field separator
							           c_proc_name           & -- procedure name
									       c_field_separator & -- field separator
										       "success"       -- message
				            severity note;
                -- error
                else
		            -- status error
                    if (v_file_status = STATUS_ERROR) then
                        assert false
			                report c_file_name                              & -- file name
							           c_field_separator                    & -- field separator
									       c_proc_name                      & -- procedure name
										       c_field_separator            & -- field separator
											       "failure : status_error"   -- message
				            severity failure;
                    -- name error 
                    elsif (v_file_status = NAME_ERROR) then
                        assert false
			                report c_file_name                              & -- file name
							           c_field_separator                    & -- field separator
									       c_proc_name                      & -- procedure name
										       c_field_separator            & -- field separator
											       "failure : name_error"     -- message
				                severity failure;
			        -- failed to open
                    else
                        assert false
			                report c_file_name                   & -- file name
 							           c_field_separator         & -- field separator 
									       c_proc_name           & -- procedure name
										       c_field_separator & -- field separator
 											       "failure"       -- message
				            severity failure;
                    end if;
		        end if;
            end procedure proc_file_rpt_open;

            -- ==========================================================================================================================================================================================
	        -- 03.01.02.02. proc_file_rpt_close
            -- ==========================================================================================================================================================================================
            procedure proc_file_rpt_close (
                 constant c_file_name : string
		        ;file     f_file      : text
            ) is 
				constant c_proc_name       : string := "proc_file_rpt_close";
			    constant c_field_separator : string := " ";			
            begin
                file_close(f_file);
		        assert false
			        report c_file_name                   & -- file name
                               c_field_separator         & -- field separator
							       c_proc_name           & -- procedure name
								       c_field_separator & -- field separator
									       "success"       -- message
			        severity note;
            end procedure proc_file_rpt_close;
	
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.03. STM
	    -- ----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
            -- ==========================================================================================================================================================================================
	        -- 03.01.02.01. proc_file_stm_open
            -- ==========================================================================================================================================================================================
            procedure proc_file_stm_open (
                 constant c_file_name : string
		        ;file     f_file      : text
            ) is                  
				constant c_proc_name       : string := "proc_file_stm_open";
			    constant c_field_separator : string := " ";
                variable v_file_status     : file_open_status;
            begin
                file_open(v_file_status,f_file,c_file_name,read_mode);
		        -- successfully opened
                if (v_file_status = OPEN_OK) then
                    assert false
			            report c_file_name                   & -- file name 
						           c_field_separator         & -- field separator
							           c_proc_name           & -- procedure name
									       c_field_separator & -- field separator
										       "success"       -- message
				            severity note;
                -- error
                else
		            -- status error
                    if (v_file_status = STATUS_ERROR) then
                        assert false
			                report c_file_name                              & -- file name
							           c_field_separator                    & -- field separator
									       c_proc_name                      & -- procedure name
										       c_field_separator            & -- field separator
											       "failure : status_error"   -- message
				            severity failure;
                    -- name error 
                    elsif (v_file_status = NAME_ERROR) then
                        assert false
			                report c_file_name                              & -- file name
							           c_field_separator                    & -- field separator
									       c_proc_name                      & -- procedure name
										       c_field_separator            & -- field separator
											       "failure : name_error"     -- message
				                severity failure;
			        -- failed to open
                    else
                        assert false
			                report c_file_name                   & -- file name
 							           c_field_separator         & -- field separator 
									       c_proc_name           & -- procedure name
										       c_field_separator & -- field separator
 											       "failure"       -- message
				            severity failure;
                    end if;
		        end if;
            end procedure proc_file_stm_open;

            -- ==========================================================================================================================================================================================
	        -- 03.01.02.02. proc_file_stm_close
            -- ==========================================================================================================================================================================================
            procedure proc_file_stm_close (
                 constant c_file_name : string
		        ;file     f_file      : text
            ) is 
				constant c_proc_name       : string := "proc_file_stm_close";
			    constant c_field_separator : string := " ";			
            begin
                file_close(f_file);
		        assert false
			        report c_file_name                   & -- file name
                               c_field_separator         & -- field separator
							       c_proc_name           & -- procedure name
								       c_field_separator & -- field separator
									       "success"       -- message
			        severity note;
            end procedure proc_file_stm_close;
	
end package body pkg_mgt_file;

-- ######################################################################################################################################################################################################
-- EOF
-- ######################################################################################################################################################################################################