-- #################################################################################################################################################################################
-- file :
--     bch_sfir_filter_4.vhd
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- objective :
--     bch_sfir_filter_4.vhd testbench file.
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- level of description :
--     behavioral
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- limitation :
--     none
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- author :
--     Tugdual LE PELLETER
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- history :
--     2024-10-19
--         file creation
-- ---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
-- table of contents :
--     01. libraries
--         01.01. standard
--         01.02. custom
--     02. entity
--     03. architecture
--         03.01. component declaration
--             03.01.01. gen_heartbeat
--             03.01.02. sfir_filter_4
--         03.02. files
--             03.02.01. LOG
--             03.02.02. RPT
--         03.03. constants
--             03.03.01. SIM
--             03.03.02. oscillator
--             03.03.03. gen_heartbeat
--             03.03.04. sfir_filter_4
--             03.03.05. arbitrary pattern generator
--             03.03.06. simulation duration
--             03.03.07. file
--         03.04. types
--             03.04.01. FSM
--                 03.04.01.01. fsm_main
--                 03.04.01.02. fsm_init
--                 03.04.01.03. fsm_test
--                 03.04.01.04. fsm_file_mgt_log
--                 03.04.01.05. fsm_file_mgt_rpt
--             03.04.02. test status
--         03.05. signals
--             03.05.01. SIM
--                 03.05.01.01. FSM
--                 03.05.01.02. files
--                 03.05.01.03. clock
--                 03.05.01.04. reset
--                 03.05.01.05. testbench
--             03.05.03. gen_heartbeat
--                 03.05.03.01. clock
--                 03.05.03.02. reset
--                 03.05.03.03. indicators
--         03.06. component instanciation
--             03.06.01. gen_heartbeat
--             03.06.02. sfir_filter_4
--         03.07. reinit
--             03.07.01. SIM
--             03.07.02. DUT    
--         03.08. clock generation
--             03.08.01. DUT
--             03.08.02. SIM
--         03.09. fsm_main
--         03.10. fsm_init
--         03.11. fsm_test
--         03.12. fsm_file_mgt_log
--         03.13. fsm_file_mgt_rpt
--         03.14. simulation abort
-- #################################################################################################################################################################################

-- #################################################################################################################################################################################
-- 01. libraries
-- #################################################################################################################################################################################
    -- =============================================================================================================================================================================
	-- 01.01. standard
    -- =============================================================================================================================================================================
    library ieee;
        use ieee.std_logic_1164.all;
	    use ieee.numeric_std.all;
	    use ieee.math_real.all;
	
    library std;
        use std.textio.all;

    -- =============================================================================================================================================================================
	-- 01.02. custom
    -- =============================================================================================================================================================================
    library work;
        use work.pkg_mgt_file.all;
		use work.pkg_gen_heartbeat.all;
	
-- #################################################################################################################################################################################
-- 02. entity
-- #################################################################################################################################################################################

entity bch_sfir_filter_4 is
end entity bch_sfir_filter_4;

-- #################################################################################################################################################################################
-- 03. architecture
-- #################################################################################################################################################################################

architecture behavioral of bch_sfir_filter_4 is

    -- =============================================================================================================================================================================
	-- 03.01. component declaration
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.01. gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component gen_heartbeat is
            generic (
	             g_clk_i_freq : integer
		        ;g_clk_o_freq : integer
	        );
            port (
	             i_clk   : in  std_logic
		        ;i_rst   : in  std_logic
		        ;o_alive : out std_logic
				;o_error : out std_logic_vector(7 downto 0)
	        );
        end component gen_heartbeat;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.01.02. sfir_filter_4
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        component sfir_filter_4 is
            generic (
        	     g_h0 : std_logic_vector(7 downto 0)
        	    ;g_h1 : std_logic_vector(7 downto 0)
        	    ;g_h2 : std_logic_vector(7 downto 0)
        	    ;g_h3 : std_logic_vector(7 downto 0)
        	);
            port (
        	     i_clk : in  std_logic
        		;i_rst : in  std_logic
        		;i_x   : in  std_logic_vector(7 downto 0)
        		;o_y   : out std_logic_vector(9 downto 0)
        	);
        end component sfir_filter_4;
        
    -- =============================================================================================================================================================================
	-- 03.02. files
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.01. LOG
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_log : text;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.02. RPT
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_rpt : text;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.02.03. STM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        file f_file_stm : text;

    -- =============================================================================================================================================================================
	-- 03.03. constants
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_sim_clk_freq      : integer := 1_000_000_000;
	    constant c_sim_clk_delay     : time    := 0.9 us;
	    constant c_sim_rst_delay     : time    := 0.3 us;
        constant c_sim_clk_period_ns : time    := integer((real(1)/real(c_sim_clk_freq))*1.0e9)*1 ns;
	    constant c_sim_clk_period    : real    := real(1)/real(c_sim_clk_freq);
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.02. oscillator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_osc_delay     : time := 2.4 us;
	    constant c_osc_freq      : integer := 100_000_000;
        constant c_osc_period_ns : time := integer((real(1)/real(c_osc_freq))*1.0e9)*1 ns;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.03. gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    constant c_dut_rst_delay    : time    := 2.5 us;
	    constant c_dut_clk_freq     : integer := c_osc_freq;
	    constant c_heartbeat_freq   : integer := 5_000_000;
		constant c_dut_clk_period   : real    := real(1)/real(c_dut_clk_freq);
	    constant c_heartbeat_period : real    := real(1)/real(c_heartbeat_freq);
	    constant c_alive_cycle_full : integer := integer(real(c_heartbeat_period)/real(c_sim_clk_period));
	    constant c_alive_cycle_half : integer := integer(real(c_alive_cycle_full)/real(2));

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.04. sfir_filter_4
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        constant c_fir_coeff_0 : std_logic_vector(7 downto 0) := "11101111";
        constant c_fir_coeff_1 : std_logic_vector(7 downto 0) := "11110101";
        constant c_fir_coeff_2 : std_logic_vector(7 downto 0) := "00011010";
        constant c_fir_coeff_3 : std_logic_vector(7 downto 0) := "00110100";
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.05. arbitrary pattern generator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_data_width       : integer := 8;
		constant c_file_stm_nb_line : integer := 2001;
	    constant c_data_freq        : integer := 100_000_000;
	    constant c_data_cnt_modulo  : integer := integer(real(c_sim_clk_freq)/real(c_data_freq));
		constant c_ratio_clk_sim_clk_dut      : integer := integer(real(c_sim_clk_freq)/real(c_dut_clk_freq));
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.06. simulation duration
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_sim_duration_factor : integer := 16;
	    constant c_sim_duration_ns     : integer := integer(real(c_sim_duration_factor)*real(c_heartbeat_period)/real(c_sim_clk_period));
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.03.07. file
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		constant c_file_log_name : string := "log_bch_sfir_filter_4_wrapper_nexys_a7_sim.csv";
		constant c_file_rpt_name : string := "rpt_bch_sfir_filter_4_wrapper_nexys_a7_sim.txt";
        constant c_file_stm_name : string := "C:\Users\Tugdual LE PELLETER\Documents\Recherche\Repositories\fir_filter_4\data\x_in_sfi_bin.txt";

	
    -- =============================================================================================================================================================================
	-- 03.04. types
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. FSM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.04.01.01. fsm_main
			-- =====================================================================================================================================================================
	        type t_fsm_main is (
	             state_fsm_main_start
                ,state_fsm_main_file_rpt_open
                ,state_fsm_main_file_log_open
                ,state_fsm_main_file_stm_open
			    ,state_fsm_main_init
		        ,state_fsm_main_run
                ,state_fsm_main_file_rpt_close
                ,state_fsm_main_file_log_close
                ,state_fsm_main_file_stm_close
		        ,state_fsm_main_stop
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.02. fsm_init
			-- =====================================================================================================================================================================
	        type t_fsm_init is (
	             state_fsm_init_idle
		        ,state_fsm_init_run
		        ,state_fsm_init_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.03. fsm_test
			-- =====================================================================================================================================================================
	        type t_fsm_test is (
	             state_fsm_test_idle
		        ,state_fsm_test_run
		        ,state_fsm_test_done
	        );
	
		    -- =====================================================================================================================================================================
			-- 03.04.01.03. fsm_test_gen_stm
			-- =====================================================================================================================================================================
	        type t_fsm_test_gen_stm is (
	             state_fsm_test_gen_stm_idle
		        ,state_fsm_test_gen_stm_run
		        ,state_fsm_test_gen_stm_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_log
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_log is (
	             state_fsm_file_mgt_log_open
				,state_fsm_file_mgt_log_write_head
	            ,state_fsm_file_mgt_log_write_data
		        ,state_fsm_file_mgt_log_close
				,state_fsm_file_mgt_log_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_rpt
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_rpt is (
	             state_fsm_file_mgt_rpt_open
	            ,state_fsm_file_mgt_rpt_write_status
		        ,state_fsm_file_mgt_rpt_close
				,state_fsm_file_mgt_rpt_done
	        );

		    -- =====================================================================================================================================================================
			-- 03.04.01.04. fsm_file_mgt_stm
			-- =====================================================================================================================================================================
	        type t_fsm_file_mgt_stm is (
	             state_fsm_file_mgt_stm_open
	            ,state_fsm_file_mgt_stm_read_data
				,state_fsm_file_mgt_stm_check_eof
		        ,state_fsm_file_mgt_stm_close
				,state_fsm_file_mgt_stm_done
	        );

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.02. test status
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	        type t_sim_test_status is (
	             TEST_OK
	            ,TEST_KO
	        );
	
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.04.01. array
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        type t_array_data is array (integer range <>) of std_logic_vector(c_data_width-1 downto 0);
	
    -- =============================================================================================================================================================================
	-- 03.05. signals
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.02. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.05.02.01. FSM
			-- =====================================================================================================================================================================
	        signal s_fsm_main_state   : t_fsm_main;
	        signal s_fsm_init_state   : t_fsm_init;
	        signal s_fsm_test_state   : t_fsm_test;
			signal s_fsm_test_gen_stm_state : t_fsm_test_gen_stm;
		    signal s_fsm_file_mgt_log : t_fsm_file_mgt_log;
		    signal s_fsm_file_mgt_rpt : t_fsm_file_mgt_rpt;
			signal s_fsm_file_mgt_stm : t_fsm_file_mgt_stm;
	
		    -- =====================================================================================================================================================================
			-- 03.05.02.02. files
			-- =====================================================================================================================================================================
		    signal s_sim_file_req_log_open  : std_logic;
		    signal s_sim_file_ack_log_open  : std_logic;
		    signal s_sim_file_req_log_close : std_logic;
		    signal s_sim_file_ack_log_close : std_logic;
		    signal s_sim_file_req_rpt_open  : std_logic;
		    signal s_sim_file_ack_rpt_open  : std_logic;
		    signal s_sim_file_req_rpt_close : std_logic;
		    signal s_sim_file_ack_rpt_close : std_logic;
		    signal s_sim_file_req_stm_open  : std_logic;
		    signal s_sim_file_ack_stm_open  : std_logic;
		    signal s_sim_file_req_stm_close : std_logic;
		    signal s_sim_file_ack_stm_close : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.03. clock
			-- =====================================================================================================================================================================
            signal s_sim_clk : std_logic;
	        signal s_osc     : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.04. reset
			-- =====================================================================================================================================================================
		    signal s_sim_rst : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.05. testbench
			-- =====================================================================================================================================================================
	        signal s_sim_cnt              : integer range 0 to c_sim_duration_ns-1;
		    signal s_sim_done             : std_logic;
		    signal s_sim_init_req         : std_logic;
		    signal s_sim_init_ack         : std_logic;
		    signal s_sim_test_req         : std_logic;
		    signal s_sim_test_ack         : std_logic;
			signal s_sim_test_ack_r       : std_logic;
			signal s_sim_test_ack_pulse   : std_logic;
			signal s_sim_test_run         : std_logic;
			signal s_sim_test_run_sr      : std_logic_vector(c_ratio_clk_sim_clk_dut-1 downto 0);
			signal s_sim_test_run_sr_tmp  : std_logic_vector(c_ratio_clk_sim_clk_dut-1 downto 0);
			signal s_sim_gen_stm          : std_logic;
		    signal s_sim_test_status      : t_sim_test_status;
			signal s_error                : std_logic;
			signal s_dut_i_data           : std_logic_vector(7 downto 0);
			
		    -- =====================================================================================================================================================================
			-- 03.05.02.05. arbitrary pattern generator
			-- =====================================================================================================================================================================
			signal s_file_stm_nb_line_cnt : integer range 0 to c_file_stm_nb_line-1;
			signal s_data                 : std_logic_vector(c_data_width-1 downto 0);
			signal s_data_array           : t_array_data(0 to c_file_stm_nb_line-1);
			signal s_data_cnt             : integer range 0 to c_data_cnt_modulo-1;
			signal s_data_idx             : integer range 0 to c_file_stm_nb_line-1;
			signal s_data_en              : std_logic;
			signal s_file_stm_eof         : std_logic;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.05.03. gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		    -- =====================================================================================================================================================================
			-- 03.05.03.01. clock
			-- =====================================================================================================================================================================
            signal s_dut_i_clk : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.03.02. reset
			-- =====================================================================================================================================================================
	        signal s_dut_i_rst : std_logic;
			signal s_dut_i_rst_n : std_logic;
			
		    -- =====================================================================================================================================================================
			-- 03.05.03.03. indicators
			-- =====================================================================================================================================================================			
		    signal s_dut_o_alive : std_logic;
			signal s_dut_o_error : std_logic_vector(7 downto 0);

begin

    -- =============================================================================================================================================================================
	-- 03.07. reset management
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_sim_rst <= '1','0' after c_sim_rst_delay;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.07.02. DUT
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        s_dut_i_rst <= '1','0' after c_dut_rst_delay;
		s_dut_i_rst_n <= not(s_dut_i_rst);

    -- =============================================================================================================================================================================
	-- 03.08. clock generation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.01. SIM
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_sim_clk : process
		begin
	        s_sim_clk <= '0';
	        wait for c_sim_clk_delay;
		    while true loop
		        s_sim_clk <= '1';
			    wait for c_sim_clk_period_ns/2;
			    s_sim_clk <= '0';
			    wait for c_sim_clk_period_ns/2;
		    end loop;
	    end process p_gen_sim_clk;

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.08.02. oscillator
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
	    p_gen_osc : process
		begin
	        s_osc <= '0';
	        wait for c_osc_delay;
		    while true loop
		        s_osc <= '1';
			    wait for c_osc_period_ns/2;
			    s_osc <= '0';
			    wait for c_osc_period_ns/2;
		    end loop;
	    end process p_gen_osc;

    -- =============================================================================================================================================================================
	-- 03.08. clock assignment
    -- =============================================================================================================================================================================
    s_dut_i_clk <= s_osc;

    -- =============================================================================================================================================================================
	-- 03.06. component instanciation
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.01. gen_heartbeat
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_dut_gen_heartbeat : gen_heartbeat
            generic map (
	             g_clk_i_freq => c_dut_clk_freq
		        ,g_clk_o_freq => c_heartbeat_freq
	        )
            port map (
	             i_clk   => s_dut_i_clk
		        ,i_rst   => s_dut_i_rst
		        ,o_alive => s_dut_o_alive
				,o_error => s_dut_o_error
	        );
			
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. s_fir_filter_4
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        inst_sfir_filter_4 : sfir_filter_4
            generic map (
                 g_h0 => c_fir_coeff_0
                ,g_h1 => c_fir_coeff_1
                ,g_h2 => c_fir_coeff_2
                ,g_h3 => c_fir_coeff_3
            )
            port map (
                 i_clk => s_dut_i_clk
        	    ,i_rst => s_dut_i_rst
        	    ,i_x   => s_dut_i_data
        	    ,o_y   => open
            );
 
    -- =============================================================================================================================================================================
	-- 03.09. fsm_main
    -- =============================================================================================================================================================================
	p_fsm_main : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_main_state <= state_fsm_main_start;
			s_sim_done <= '0';
			s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
			s_sim_file_req_stm_open <= '0';
			s_sim_file_req_stm_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_done <= '0';
            s_sim_init_req <= '0';
			s_sim_test_req <= '0';
			s_sim_file_req_log_open <= '0';
			s_sim_file_req_log_close <= '0';
			s_sim_file_req_rpt_open <= '0';
			s_sim_file_req_rpt_close <= '0';
			s_sim_file_req_stm_open <= '0';
			s_sim_file_req_stm_close <= '0';
		    case s_fsm_main_state is
			    -- wait for DUT reset deassertion
				when state_fsm_main_start =>
				    if (s_dut_i_rst = '0') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_open;
						s_sim_file_req_rpt_open <= '1';
					end if;
				-- wait for RPT file to be opened
			    when state_fsm_main_file_rpt_open =>
				    if (s_sim_file_ack_rpt_open = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_open;
					    s_sim_file_req_log_open <= '1';
					end if;
				-- wait for LOG file to be opened
				when state_fsm_main_file_log_open =>
				    if (s_sim_file_ack_log_open = '1') then
					    s_fsm_main_state <= state_fsm_main_file_stm_open;
						s_sim_file_req_stm_open <= '1';
					end if;
				-- wait for STM file to be opened
				when state_fsm_main_file_stm_open =>
				    if (s_sim_file_ack_stm_open = '1') then
					    s_fsm_main_state <= state_fsm_main_init;
						s_sim_init_req <= '1';
					end if;
				-- waiting for init done
				when state_fsm_main_init =>
				    if (s_sim_init_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_run;
					    s_sim_test_req <= '1';
					end if;
				-- waiting for test done
				when state_fsm_main_run =>
                    if (s_sim_test_ack = '1') then
					    s_fsm_main_state <= state_fsm_main_file_log_close;
						s_sim_file_req_log_close <= '1';
					end if;
				-- waiting for data file to be closed
				when state_fsm_main_file_log_close =>
                    if (s_sim_file_ack_log_close = '1') then
					    s_fsm_main_state <= state_fsm_main_file_rpt_close;
						s_sim_file_req_rpt_close <= '1';
					end if;
				-- waiting for SIM report file to be closed
				when state_fsm_main_file_rpt_close =>
                    if (s_sim_file_ack_rpt_close = '1') then
					    s_fsm_main_state <= state_fsm_main_file_stm_close;
				        s_sim_file_req_stm_close <= '1';
					end if;
				-- waiting for SIM report file to be closed
				when state_fsm_main_file_stm_close =>
                    if (s_sim_file_ack_stm_close = '1') then
					    s_fsm_main_state <= state_fsm_main_stop;
				        s_sim_done <= '1';
					end if;
				-- test stopped
                when state_fsm_main_stop =>
                    null;
			end case;
		end if;
	end process p_fsm_main;

    -- =============================================================================================================================================================================
	-- 03.10. fsm_init
    -- =============================================================================================================================================================================
	fsm_init : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_init_state <= state_fsm_init_idle;
			s_sim_init_ack <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_init_ack <= '0';
		    case s_fsm_init_state is
			    -- waiting for init request
			    when state_fsm_init_idle =>
				    if (s_sim_init_req = '1') then
					    s_fsm_init_state <= state_fsm_init_run;
					end if;
				-- running init
				when state_fsm_init_run =>
					s_fsm_init_state <= state_fsm_init_done;
                    s_sim_init_ack <= '1';
				-- init done
                when state_fsm_init_done =>
				    null;
			end case;
		end if;
	end process fsm_init;

    -- =============================================================================================================================================================================
	-- 03.11. fsm_test
    -- =============================================================================================================================================================================
	p_fsm_test : process(s_sim_rst,s_sim_clk)
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_test_state <= state_fsm_test_idle;
			s_sim_test_run <= '0';
			s_sim_test_status <= TEST_OK;
		elsif (rising_edge(s_sim_clk)) then
			s_sim_test_run <= '0';
		    case s_fsm_test_state is
			    -- waiting for test request
			    when state_fsm_test_idle =>
				    if (s_sim_test_req = '1') then
					    s_sim_test_run <= '1';
					    s_fsm_test_state <= state_fsm_test_run;
					end if;
				-- running test
				when state_fsm_test_run =>
					-- parsing data vector
					if (s_sim_test_ack_pulse = '1') then
					    s_fsm_test_state <= state_fsm_test_done;
						s_sim_test_status <= TEST_OK;
					end if;
				-- test done
                when state_fsm_test_done =>
                    null;
			end case;
		end if;
	end process p_fsm_test;

    -- =============================================================================================================================================================================
	-- 03.12. stimuli generator
    -- =============================================================================================================================================================================
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. Regenerate request pulse (From fast to slow clock domain)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        p_sim_test_run_sr : process(s_sim_rst,s_sim_clk)
		begin
		    if (s_sim_rst = '1') then
			    s_sim_test_run_sr <= (others => '0');
			elsif (rising_edge(s_sim_clk)) then
			    s_sim_test_run_sr <= s_sim_test_run_sr(s_sim_test_run_sr'high-1 downto 0) & s_sim_test_run;
			end if;
		end process p_sim_test_run_sr;
 
        s_sim_test_run_sr_tmp(0) <= s_sim_test_run_sr(0);
		
		or_gen_test_run : for i in 1 to c_ratio_clk_sim_clk_dut-1 generate
		    s_sim_test_run_sr_tmp(i) <= s_sim_test_run_sr(i) or s_sim_test_run_sr_tmp(i-1);
		end generate or_gen_test_run;
		
		s_sim_gen_stm <= s_sim_test_run_sr_tmp(s_sim_test_run_sr_tmp'length-1);

	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
		-- 03.06.02. Generate stimuli (DUT clock domain)
	    -- -------------------------------------------------------------------------------------------------------------------------------------------------------------------------
        p_fsm_test_gen_stm : process(s_dut_i_rst,s_dut_i_clk)
	    begin
	        if (s_dut_i_rst = '1') then
			    s_fsm_test_gen_stm_state <= state_fsm_test_gen_stm_idle;
				s_data_idx <= 0;
				s_dut_i_data <= (others => '0');
				s_sim_test_ack <= '0';
	    	elsif (rising_edge(s_dut_i_clk)) then
			    s_sim_test_ack <= '0';
                case s_fsm_test_gen_stm_state is
				     when state_fsm_test_gen_stm_idle =>
					    if (s_sim_gen_stm = '1') then
						    s_fsm_test_gen_stm_state <= state_fsm_test_gen_stm_run;
						end if;
				    -- parsing stimuli vector
					 when state_fsm_test_gen_stm_run =>
					    -- feeding filter with data
					    s_dut_i_data <= s_data_array(s_data_idx);
					    if (s_data_idx = c_file_stm_nb_line-1) then
						   s_data_idx <= 0;
						   s_sim_test_ack <= '1';
						   s_fsm_test_gen_stm_state <= state_fsm_test_gen_stm_done;
						else
						   s_data_idx <= s_data_idx + 1;
						end if;
					 when state_fsm_test_gen_stm_done =>
					    null;
				end case;
	    	end if;
	    end process p_fsm_test_gen_stm;

        p_test_ack_pulse : process(s_sim_rst,s_sim_clk)
		begin
		    if (s_sim_rst = '1') then
			    s_sim_test_ack_r <= '0';
				s_sim_test_ack_pulse <= '0';
			elsif (rising_edge(s_sim_clk)) then
			    if (s_sim_test_ack_r = '0' and s_sim_test_ack_r = '1') then
				    s_sim_test_ack_pulse <= '1';
				else
				    s_sim_test_ack_pulse <= '0';
				end if;
			end if;
		end process p_test_ack_pulse;

    -- =============================================================================================================================================================================
	-- 03.12. fsm_file_mgt_stm
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_stm : process(s_sim_rst,s_sim_clk)
		constant c_justified  : side   := right;
		constant c_field      : width  := 0;
		constant c_unit       : time   := ns;
		constant c_separator  : string := ",";
		constant c_value_head : string := "time,data";
	    variable v_value_time : time;
		variable v_value_data : bit_vector(c_data_width-1 downto 0);
		variable v_value_foot : string(1 to 7);
		variable v_line       : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_stm <= state_fsm_file_mgt_stm_open;
		    s_sim_file_ack_stm_open <= '0';
			s_sim_file_ack_stm_close <= '0';
			s_file_stm_nb_line_cnt <= 0;
			s_data_array <= (others => (others => '0'));
			s_file_stm_eof <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_stm_open <= '0';
			s_sim_file_ack_stm_close <= '0';
            case s_fsm_file_mgt_stm is
                -- open file
			    when state_fsm_file_mgt_stm_open =>
				    if (s_sim_file_req_stm_open = '1') then
					    s_fsm_file_mgt_stm <= state_fsm_file_mgt_stm_read_data;
						s_sim_file_ack_stm_open <= '1';
						proc_file_stm_open(c_file_stm_name,f_file_stm);
					end if;
				-- read data from file (at least one line)
				when state_fsm_file_mgt_stm_read_data =>
                    readline(f_file_stm,v_line);
                    read(v_line,v_value_data);
					s_data_array(s_file_stm_nb_line_cnt) <= to_stdlogicvector(v_value_data);
                    s_fsm_file_mgt_stm <= state_fsm_file_mgt_stm_check_eof;
                -- close file
				when state_fsm_file_mgt_stm_check_eof =>
				    if (s_file_stm_nb_line_cnt = c_file_stm_nb_line-1) then
					    s_file_stm_nb_line_cnt <= 0;
						s_file_stm_eof <= '1';
					    s_fsm_file_mgt_stm <= state_fsm_file_mgt_stm_close;
					else
					    s_file_stm_nb_line_cnt <= s_file_stm_nb_line_cnt + 1;
					    s_fsm_file_mgt_stm <= state_fsm_file_mgt_stm_read_data;
					end if;
				when state_fsm_file_mgt_stm_close =>
				    if (s_sim_file_req_stm_close = '1') then
					    s_fsm_file_mgt_stm <= state_fsm_file_mgt_stm_done;
				        s_sim_file_ack_stm_close <= '1';
                        proc_file_stm_close(c_file_stm_name,f_file_stm);
					end if;
				-- done
				when state_fsm_file_mgt_stm_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_stm;

    -- =============================================================================================================================================================================
	-- 03.12. fsm_file_mgt_log
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_log : process(s_sim_rst,s_sim_clk)
		constant c_justified  : side   := right;
		constant c_field      : width  := 0;
		constant c_unit       : time   := ns;
		constant c_separator  : string := ",";
		constant c_value_head : string := "time,data";
	    variable v_value_time : time;
		variable v_value_data : string(1 to 4);
		variable v_value_foot : string(1 to 7);
		variable v_line       : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_open;
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_log_open <= '0';
			s_sim_file_ack_log_close <= '0';
            case s_fsm_file_mgt_log is
                -- open file
			    when state_fsm_file_mgt_log_open =>
				    if (s_sim_file_req_log_open = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_head;
						s_sim_file_ack_log_open <= '1';
						proc_file_log_open(c_file_log_name,f_file_log);
					end if;
				-- write header
				when state_fsm_file_mgt_log_write_head =>
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_write_data;
						write(v_line,c_value_head,c_justified,c_field);
	                    writeline(f_file_log,v_line);
				-- write data
				when state_fsm_file_mgt_log_write_data =>
				    if (s_sim_file_req_log_close = '1') then
					    s_fsm_file_mgt_log <= state_fsm_file_mgt_log_close;
						-- timestamp
						v_value_time := now;
						write(v_line,v_value_time,c_justified,c_field,c_unit);
						-- separator
						write(v_line,c_separator,c_justified,c_field);
						-- data value
						v_value_data := "NONE";
					    write(v_line,v_value_data,c_justified,c_field);
	                    writeline(f_file_log,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_log_close =>
					s_fsm_file_mgt_log <= state_fsm_file_mgt_log_done;
				    s_sim_file_ack_log_close <= '1';
                    proc_file_log_close(c_file_log_name,f_file_log);
				-- done
				when state_fsm_file_mgt_log_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_log;

    -- =============================================================================================================================================================================
	-- 03.13. fsm_file_mgt_rpt
    -- =============================================================================================================================================================================
	p_fsm_file_mgt_rpt : process(s_sim_rst,s_sim_clk)
		constant c_justified    : side  := right;
		constant c_field        : width := 0;
		variable v_value_status : string(1 to 7);
		variable v_line         : line;
	begin
	    if (s_sim_rst = '1') then
		    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_open;
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
		elsif (rising_edge(s_sim_clk)) then
		    s_sim_file_ack_rpt_open <= '0';
			s_sim_file_ack_rpt_close <= '0';
            case s_fsm_file_mgt_rpt is
                -- open file
			    when state_fsm_file_mgt_rpt_open =>
				    if (s_sim_file_req_rpt_open = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_write_status;
						s_sim_file_ack_rpt_open <= '1';
						proc_file_rpt_open(c_file_rpt_name,f_file_rpt);
					end if;
				-- write status
				when state_fsm_file_mgt_rpt_write_status =>
				    if (s_sim_file_req_rpt_close = '1') then
					    s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_close;
					    -- write test status
					    case s_sim_test_status is
					        when TEST_OK => v_value_status := "TEST_OK";
						    when others  => v_value_status := "TEST_KO";
					    end case;
					    write(v_line,v_value_status,c_justified,c_field);
	                    writeline(f_file_rpt,v_line);
					end if;
                -- close file
				when state_fsm_file_mgt_rpt_close =>
					s_fsm_file_mgt_rpt <= state_fsm_file_mgt_rpt_done;
				    s_sim_file_ack_rpt_close <= '1';
                    proc_file_rpt_close(c_file_rpt_name,f_file_rpt);
				-- done
				when state_fsm_file_mgt_rpt_done  =>
				    null;
			end case;
		end if;
	end process p_fsm_file_mgt_rpt;

    -- =============================================================================================================================================================================
	-- 03.14. error detection
    -- =============================================================================================================================================================================
	p_check_dut_error : process(s_dut_i_rst,s_sim_clk)
	    variable v_error : std_logic;
	begin
	    if (s_dut_i_rst = '1') then
	        v_error := '0';
			s_error <= '0';
	    elsif (rising_edge(s_sim_clk)) then
		    v_error := '0';
			-- parsing error vector
		    for i in 0 to s_dut_o_error'length-1 loop
		        -- error detected
			    if (s_dut_o_error(i) = '1') then
				    v_error := '1';
				end if;
			end loop;
			s_error <= v_error;
		end if;
	end process p_check_dut_error;	
	
    -- =============================================================================================================================================================================
	-- 03.14. simulation abort : clock ratio error
    -- =============================================================================================================================================================================
	p_sim_abort : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_error = '1') then
			    assert false 
				    report "end of simulation - DUT error detected" 
					    severity failure;
			end if;
		end if;
	end process p_sim_abort;

    -- =============================================================================================================================================================================
	-- 03.14. end of simulation
    -- =============================================================================================================================================================================
	p_sim_end : process(s_sim_clk)
	begin
		if (rising_edge(s_sim_clk)) then
            if (s_sim_done = '1') then
			    assert false 
				    report "end of simulation - success" 
					    severity failure;
			end if;
		end if;
	end process p_sim_end;

end architecture behavioral;

-- #################################################################################################################################################################################
-- EOF
-- #################################################################################################################################################################################